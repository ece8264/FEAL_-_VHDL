library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity reg128 is
	port(   CLK,RST,EN_INPUT: in std_logic;
		DATA_IN: in std_logic_vector(127 downto 0);
		DATA_OUT: out std_logic_vector(127 downto 0));
	
end reg128;

architecture my_arch of reg128 is

signal RegVal: std_logic_vector(127 downto 0);

begin
	
process(RST,CLK)

variable  RegVal: std_logic_vector(127 downto 0);

begin 

if(RST = '1') then 
RegVal := (others => '0');
DATA_OUT <= RegVal;
elsif (CLK'event AND CLK = '1') then
	if(EN_INPUT = '1') then 
	RegVal := DATA_IN;
	DATA_OUT <= RegVal;
	end if;
end if;
end process;

end my_arch;
