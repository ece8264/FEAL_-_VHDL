library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity MUX96_32 is
	port(   X0 : in std_logic_vector(31 downto 0);
	  	X1 : in std_logic_vector(31 downto 0);
		X2 : in std_logic_vector(31 downto 0);
		MUX96_32_OUT : out std_logic_vector(31 downto 0);
		SEL: in integer range 0 to 2 );
end MUX96_32;


architecture myarch of MUX96_32 is
begin 
with SEL select MUX96_32_OUT <= 
	X0 when 0,
	X1 when 1,
	X2 when others;
	   
end myarch;
	